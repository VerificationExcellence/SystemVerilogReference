//---------------------
// Monitor class
//---------------------
class eth_packet_mon_c;

 //Virtual interface to sample signals
 //TBD


 //Method to sample signal on a port and then
 //create a packet class and print it

endclass
