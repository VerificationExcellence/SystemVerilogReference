bit  a, b, c, d, e; 
always @(a, b, c) begin
  e =  a & b & c &d 
end
