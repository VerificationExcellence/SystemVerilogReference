//----------------
//Packet driver class
//----------------
class eth_packet_drv_c;

  //Use a virtual interface that points to same interface

  //Use a mailbox to receive packets from generator

  //Implement a function that can drive the design interface signals
  //as per the packet fields

endclass
