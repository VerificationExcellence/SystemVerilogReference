//---------------------
// Monitor class
//---------------------
class eth_packet_mon_c;

 //Virtual interface to sample signals
 //TBD


 //Method to sample signal on a port and then
 //create a packet class and print it

 //Use a mailbox to put the packets monitored on both input
 // and output ports

endclass
