interface  rr_assert_if(
  input logic reset,
  input logic clk,
  input logic[3:0] req,
  input logic[3:0] grant
);
  
  
  
endinterface
