//------------------------------------
// This will be a stand alone module that illustrates usages of several of
// SV basic data types and usages
// This can be compiled as a stand alone file
// Students can experiment  by compiling and simulating this file
// and observing the behavior
//------------------------------------
module data_types_eg;


//bit vs logic difference
//packed vs unpacked



endmodule
