//-----------------------------
//Packet generator class
//-----------------------------
class eth_packet_gen_c;

  //Implement a random member for number of packets to be generated

  //Implement a method which when called should create so many packets - after randomizing each

  //Use a mail box and put these generated packets into that
  //This mailbox will be later used by the driver

  //TBD

endclass
